module moduleName #(
    parameters
) (
    ports
);
    
endmodul